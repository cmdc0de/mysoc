module soc
begin
endmodule
